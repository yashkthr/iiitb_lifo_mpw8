// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq
);
  

    wire [`MPRJ_IO_PADS-1:0] io_in;
    wire [`MPRJ_IO_PADS-1:0] io_out;
    wire [`MPRJ_IO_PADS-1:0] io_oeb;



    // IO
    assign clk = wb_clk_i;
    assign Rst = wb_rst_i;
    assign {dataIn,RW,EN} = io_in[37:32];
    assign io_out[37:32] = {dataOut,EMPTY,FULL};
    assign io_oeb = 0;

    // IRQ
    assign irq = 3'b000;	// Unused

    
    wire dataIn;
    wire dataOut; 
    wire RW; 
    wire EN;
    wire Rst;
    wire EMPTY;
    wire FULL;
    wire clk;

    iiitb_lifo i1 (dataIn, dataOut, RW, EN,
                   Rst,
                   EMPTY,
                   FULL,
                   clk);

endmodule

module iiitb_lifo( dataIn, dataOut, RW, EN,
                   Rst,
                   EMPTY,
                   FULL,
                   clk
                  );
input [3:0]  dataIn;
input        RW,
             EN,
             Rst,
             clk;
     
output  reg EMPTY,
            FULL;    
output reg [3:0] dataOut;
reg [3:0] stack_mem[0:3];
reg  [2:0] SP;
integer i;
  always @ (posedge clk)
begin
 if (EN==0);
 else begin
    if (Rst==1) begin
      SP       = 3'd4;
      EMPTY    = SP[2];
      dataOut  = 4'h0;
      for (i=0;i<4;i=i+1) begin
        stack_mem[i]= 0;
      end
     end
  else if (Rst==0) begin
    FULL = SP? 0:1;
    EMPTY  = SP[2];
    dataOut = 4'hx;
    if (FULL == 1'b0 && RW == 1'b0) begin
       SP            = SP-1'b1;
       FULL          = SP? 0:1;
       EMPTY         = SP[2];
       stack_mem[SP] = dataIn;
     end
   else if (EMPTY == 1'b0 && RW == 1'b1) begin
       dataOut  = stack_mem[SP];
       stack_mem[SP] = 0;
       SP  = SP+1;
       FULL  = SP? 0:1;
       EMPTY  = SP[2];
    end
   else;
  end
  else;
 end
end
endmodule
`default_nettype wire
